// Module Name:     sram
// Author:          WuHan University  clong
// Date Created:    1-June-2020


package apb_global_pkg;
    // include global defines
    `include "tb_defines.sv"

endpackage